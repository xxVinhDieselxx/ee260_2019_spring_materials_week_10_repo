module problem_3(clk, x, y);
  input clk;
  input x;
  output reg y;
  /* your code */
endmodule