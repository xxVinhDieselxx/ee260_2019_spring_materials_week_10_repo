`timescale 1 ns / 100 ps
module problem_7_tb();
  /* your code */
endmodule
